* TLC2254 OPERATIONAL AMPLIFIER "MACROMODEL" SUBCIRCUIT
* CREATED USING PARTS RELEASE 4.03 ON 11/07/94 AT 09:12
* (5V MODEL)
* CONNECTIONS:   NON-INVERTING INPUT
*                | INVERTING INPUT
*                | | POSITIVE POWER SUPPLY
*                | | | NEGATIVE POWER SUPPLY
*                | | | | OUTPUT
*                | | | | |
.SUBCKT TLC2254  1 2 3 4 5
*
  C1   11 12 6.369E-12
  C2    6  7 25.00E-12
  CSS  10 99 3.182E-12
  DC    5 53 DX
  DE   54  5 DX
  DLP  90 91 DX
  DLN  92 90 DX
  DP    4  3 DX
  EGND 99  0 POLY(2) (3,0) (4,0) 0 .5 .5
  FB    7 99 POLY(5) VB VC VE VLP VLN 0 57.62E6 -60E6 60E6 60E6 -60E6
  GA    6  0 11 12 26.86E-6
  GCM   0  6 10 99 2.686E-9
  ISS   3 10 DC 3.100E-6
  HLIM 90  0 VLIM 1K
  J1   11  2 10 JX
  J2   12  1 10 JX
  R2    6  9 100.0E3
  RD1 60 11 37.23E3
  RD2 60 12 37.23E3
  RO1   8  5 84
  RO2   7 99 84
  RP    3  4 71.43E3
  RSS  10 99 64.52E6
  VAD  60 4 -.5
  VB    9  0 DC 0
  VC 3 53 DC .605
  VE   54  4 DC .605
  VLIM  7  8 DC 0
  VLP  91  0 DC -.235
  VLN 0 92 DC 7.500
.MODEL DX D(IS=800.0E-18)
.MODEL JX PJF(IS=500.0E-15 BETA=139E-6 VTO=-.05)
.ENDS
